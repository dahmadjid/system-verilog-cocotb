module ent (
    input  logic a,
    output logic b
);
  always_comb begin
    b = a;
  end
endmodule
